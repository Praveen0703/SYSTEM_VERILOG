module onedimensional_array;
  int array[2];
  initial begin
    foreach(array[i])begin
      array[i]=$random;
    end
    $display("output=%p",array);
  end
endmodule
output='{303379748, -1064739199}

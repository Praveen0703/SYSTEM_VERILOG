module threedimensional_array;
  int array[2:0][3:0][4:0];
  initial begin
    foreach(array[i,k,l])begin
      array[i][k][l]=$random;
    end
    $display("array=%p",array);
  end
endmodule
      array='{'{'{303379748, -1064739199, -2071669239, -1309649309, 112818957}, '{1189058957, -1295874971, -1992863214, 15983361, 114806029}, '{992211318, 512609597, 1993627629, 1177417612, 2097015289}, '{-482925370, -487095099, -720121174, 1924134885, -1143836041}}, '{'{-1993157102, 1206705039, 2033215986, -411658546, -201295128}, '{-490058043, 777537884, -561108803, -1767155667, -1297668507}, '{-1309711773, 91457290, -1069866368, 274997536, 1433945514}, '{-825439075, -887079274, -1987856365, -2034485235, -1448618413}}, '{'{899669355, -358208811, -2129180158, -682213714, 251652381}, '{-406490417, 293882147, 84501770, -445445430, -1640936388}, '{2036907506, 1160667530, 549761857, -330615592, 1008792440}, '{-997584247, 1975848427, 1526883766, 1665923526, 1460999086}}}
